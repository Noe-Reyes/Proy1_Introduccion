module and_gate
(
    input a,
    input b,
    output y
);
    assign y = a & b;
    // Aun no le entiendo al pinche programa.
    //Creo que al menos lo mas facil ya lo se hacer.
    // Vamos a probar otra modificacion, para saber como funciona.
    // Asi se hace un cambio.
endmodule